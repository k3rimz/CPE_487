--start
--library declarations
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY accelerometer IS
    PORT (

    );
END  accelerometer;

  
  
ARCHITECTURE Behavioral OF  accelerometer IS

END Behavioral;
